// module control (
//     // IN
//     input logic [6:0] op,
//     input logic [2:0] func3,
//     input logic [6:0] func7,
//     input logic alu_zero,

//     // OUT
//     output logic [2:0] alu_control,
//     output logic [1:0] imm_source,
//     output logic mem_write,
//     output logic reg_write
// );

// /**
// * MAIN DECODER
// */

// always_comb begin

//         // --- 1. DECODE LOGIC ---
//         if (op == 7'b0000011) begin : LW_DECODE
//             // I-type (lw)
//             reg_write   = 1'b1;
//             imm_source  = 2'b00;
//             mem_write   = 1'b0;
//             alu_control = 3'b000; // ADD
//         end 
//         else if (op == 7'b0100011) begin : SW_DECODE
//             // S-type (sw)
//             reg_write   = 1'b0;
//             imm_source  = 2'b01;
//             mem_write   = 1'b1;
//             alu_control = 3'b000; // ADD
//         end
//         else begin : DEFAULT_DECODE
//             // This is your "Everything Else" catch-all
//             reg_write   = 1'b0;
//             mem_write   = 1'b0;
//             imm_source  = 2'b00;
//             alu_control = 3'b111;
//         end
// end
    
// endmodule



module control (
    // IN
    input logic [6:0] op,
    input logic [2:0] func3,
    input logic [6:0] func7,
    input logic alu_zero,

    // OUT
    output logic [2:0] alu_control,
    output logic [1:0] imm_source,
    output logic mem_write,
    output logic reg_write
);

/**
* MAIN DECODER
*/

logic [1:0] alu_op;
always_comb begin
    case (op)
        // I-type (lw)
        7'b0000011 : begin
            reg_write = 1'b1;
            imm_source = 2'b00;
            mem_write = 1'b0;
            alu_op = 2'b00;
        end
        // S-Type (sw)
        7'b0100011 : begin
            reg_write = 1'b0;
            imm_source = 2'b01;
            mem_write = 1'b1;
            alu_op = 2'b00;
        end
        // EVERYTHING ELSE
        default: begin
            reg_write = 1'b0;
            imm_source = 2'b00;
            mem_write = 1'b0;
            alu_op = 2'b00;
        end
    endcase
end

/**
* ALU DECODER
*/

always_comb begin
    case (alu_op)
        // LW, SW
        2'b00 : alu_control = 3'b000;
        // EVERYTHING ELSE
        default: alu_control = 3'b111;
    endcase
end
    
endmodule